// ============================================================================
//        __
//   \\__/ o\    (C) 2021  Robert Finch, Waterloo
//    \  __ /    All rights reserved.
//     \/_//     robfinch<remove>@finitron.ca
//       ||
//
//	Thor2021_hiAmt.sv
//  - head pointers increment amount
//
//
// BSD 3-Clause License
// Redistribution and use in source and binary forms, with or without
// modification, are permitted provided that the following conditions are met:
//
// 1. Redistributions of source code must retain the above copyright notice, this
//    list of conditions and the following disclaimer.
//
// 2. Redistributions in binary form must reproduce the above copyright notice,
//    this list of conditions and the following disclaimer in the documentation
//    and/or other materials provided with the distribution.
//
// 3. Neither the name of the copyright holder nor the names of its
//    contributors may be used to endorse or promote products derived from
//    this software without specific prior written permission.
//
// THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS"
// AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE
// IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE
// DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTORS BE LIABLE
// FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL
// DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR
// SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER
// CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY,
// OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE
// OF THIS SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
//                                                                          
// ============================================================================

import Thor2021_pkg::*;

module Thor2021_hiAmt(rob, commit0_v, commit1_v, heads, tails, amt_o);
parameter RENTRIES = `RENTRIES;
input sReorderEntry rob [0:RENTRIES-1];
input commit0_v;
input commit1_v;
input SrcId heads [0:RENTRIES-1];
input SrcId tails [0:1];
output reg [2:0] amt_o;

reg [2:0] amt;
SrcId nxtrb;

// Determine amount to advance reorder head pointer by. Based on number of
// consecutive valid commits. Also up to four additional slot that have been
// marked invalid may be advanced past.
always_comb
begin
	if (commit0_v & commit1_v)
		amt = 3'd2;
	else if (commit0_v)
		amt = 3'd1;
	else
		amt = 3'd0;

	// Now search ahead for invalid entries that can be skipped over.
	nxtrb = (heads[0] + amt) % RENTRIES;
	if (rob[nxtrb].state==RS_INVALID && heads[nxtrb]!=tails[0]) begin
		amt = amt + 4'd1;
		nxtrb = (heads[0] + amt) % RENTRIES;
		if (rob[nxtrb].state==RS_INVALID && heads[nxtrb]!=tails[0]) begin
			amt = amt + 4'd1;
			nxtrb = (heads[0] + amt) % RENTRIES;
			if (rob[nxtrb].state==RS_INVALID && heads[nxtrb]!=tails[0]) begin
				amt = amt + 4'd1;
				nxtrb = (heads[0] + amt) % RENTRIES;
				if (rob[nxtrb].state==RS_INVALID && heads[nxtrb]!=tails[0]) begin
					amt = amt + 4'd1;
					nxtrb = (heads[0] + amt) % RENTRIES;
				end
			end
		end
	end
	amt_o = amt;
end

endmodule
