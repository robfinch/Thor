module Thor2022_gpr_file();
endmodule